module top(
        input a,
        output b
        
);

        always @(*)
        begin
                b = a;
        end

endmodule
